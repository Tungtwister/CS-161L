`timescale 1ns / 1ps

`define FP_SIZE 32

module FP_Adder(
input clk,
input rst,
input enable,
output reg valid,
input [31:0] A,
input [31:0] B,
output reg[`FP_SIZE-1:0] result
);
// Implement your code here
//Combinational Part
reg [31:0] yourresult;
reg [31:0] C;
reg signA, signB; //sign bits for A and B
reg givenSA, givenSB; //given sign bits for A and B
reg signC;
reg [7:0] expA, expB; //exponent bits for A and B
reg [7:0] expC;
reg [22:0] mantisA, mantisB; //mantissa bits for A and B
reg [23:0] exManA, exManB; //extended mantissa A and B
reg [32:0] tmp;
reg tmpS;
reg [7:0] tmpE;
reg [23:0] tmpM;
integer tmpI;
integer expDif;
reg carryout = 0;
reg [23:0] mantisC;
reg [7:0] shift;
integer i = 0;

always @ (*) begin
//step 1
signA = A[31]; //Separate sign bit from inputs A and B
signB = B[31];
givenSA = A[31]; //Separate sign bit from inputs A and B
givenSB = B[31];

expA = A[30:23]; //Separate exponent bits from inputs A and B
expB = B[30:23];

mantisA = A[22:0]; //Separate mantissa bits from inputs A and B
mantisB = B[22:0];
//--------------------------------------------------------------
exManA = {{1'b1},{mantisA}};
exManB = {{1'b1},{mantisB}};
//$display("%b",signB);
//$display("%b",expB);
//$display("%b",exManB);

//step 2
if(expB > expA)
begin
	tmpS = signA;
	tmpE = expA;
	tmpM = exManA;
	signA = signB;
	expA = expB;
	exManA = exManB;
	signB = tmpS;
	expB = tmpE;
	exManB = tmpM;
end
	expDif = expA - expB; //exponent difference
//step 3
exManB = exManB >> expDif;
//step 4
if(signA != signB)
begin
tmp = {{signB},{expB},{exManB}};
tmp = -tmp;
signB = tmp[32];
expB = tmp[31:24];
exManB = tmp[23:0];
end
//step 5
{carryout, mantisC} = exManA + exManB;
//step 6
if(givenSA != givenSB)
begin
	{carryout, mantisC} = -{carryout, mantisC};
end
//step 7
shift = 0;
if((givenSA == givenSB) && (carryout == 1'b1))
begin
	mantisC = mantisC >> 1;
	mantisC[23] = 1'b1;
	shift = 1;
end
else
begin
	for(i =0; i<24; i=i+1)
	begin
			if(mantisC[23] == 0)
			begin
			mantisC = mantisC << 1;
			shift = shift + 1;
			end
	end
end

//step 8
if((givenSA != givenSB) && (B[30:0] > A[30:0]))
begin
signC = givenSB;
expC = expB + 1;
end
else
begin
signC = givenSA;
expC = expA + shift;
end
//step 9

if(shift == 24)
begin
C = 32'h0;
end
else
begin
C = {{signC},{expC},{mantisC[22:0]}};
end

yourresult = C;
end

// Sequential Part
always @(posedge clk) begin
if (rst) begin
result <= 0;
valid <= 0;
end
else begin
result <= yourresult;
valid <= enable;
end
end
endmodule
